----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:45:44 07/06/2016 
-- Design Name: 
-- Module Name:    MUL2_COM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUL2_COM is
    Port ( I : in  STD_LOGIC_VECTOR (1 downto 0);
           S : in  BIT;
           Y : out  STD_LOGIC);
end MUL2_COM;

architecture Behavioral of MUL2_COM is

begin
Y <= I(0) when S='0' else
	  I(1);

end Behavioral;

