--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   19:19:36 07/06/2016
-- Design Name:   
-- Module Name:   E:/VHDL/fzyserial4/fzyserial4_tb.vhd
-- Project Name:  fzyserial4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: fzyserial4
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY fzyserial4_tb IS
END fzyserial4_tb;
 
ARCHITECTURE behavior OF fzyserial4_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT fzyserial4
    PORT(
         A : IN  std_logic;
         clk : IN  std_logic;
         B : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic := '0';
   signal clk : std_logic := '0';

 	--Outputs
   signal B : std_logic:= '0';

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: fzyserial4 PORT MAP (
          A => A,
          clk => clk,
          B => B
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for clk_period;	
		A <='1';
		wait for clk_period;
		A <='0';
		wait for clk_period;
		A <='1';
		wait for clk_period;	
		A <='0';
		wait for clk_period;
		A <='1';
		wait for clk_period;
		A <='0';
		wait for clk_period;
		A <='1';
		wait for clk_period;
		A <='0';
	

      wait;
   end process;

END;
